`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:54:33 05/07/2016 
// Design Name: 
// Module Name:    Select_Wd 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Select_Wd(
input WrRegData,
input [31:0] in0,
input [31:0] in1,
output [31:0] out
    );
	always @ (*)
		

endmodule
